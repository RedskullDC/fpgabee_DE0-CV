library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;


entity pcu_rom is
	port
	(
		clock : in std_logic;
		clken : in std_logic;
		addr : in std_logic_vector(11 downto 0);
		dout : out std_logic_vector(7 downto 0)
	);
end pcu_rom;
 
architecture behavior of pcu_rom is 
	type mem_type is array(0 to 4095) of std_logic_vector(7 downto 0);	signal rom : mem_type := 
	(
	x"c3", x"02", x"0a", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"c3", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"ed", x"73", x"b2", x"42", x"31", x"c2", x"42", x"f5", x"c5", x"d5", x"e5", x"dd", x"e5", x"fd", x"e5", x"ed", 
	x"7b", x"b4", x"42", x"fd", x"e1", x"dd", x"e1", x"e1", x"d1", x"c1", x"f1", x"c9", x"f5", x"c5", x"d5", x"e5", 
	x"dd", x"e5", x"fd", x"e5", x"ed", x"73", x"b4", x"42", x"31", x"b6", x"42", x"fd", x"e1", x"dd", x"e1", x"e1", 
	x"d1", x"c1", x"f1", x"ed", x"7b", x"b2", x"42", x"d3", x"80", x"ed", x"45", x"e5", x"d5", x"db", x"82", x"5f", 
	x"db", x"83", x"cb", x"7f", x"20", x"05", x"cd", x"1c", x"01", x"18", x"f2", x"16", x"00", x"21", x"68", x"03", 
	x"19", x"19", x"cb", x"47", x"28", x"01", x"23", x"7e", x"fe", x"1c", x"20", x"08", x"db", x"81", x"ee", x"03", 
	x"d3", x"81", x"18", x"d9", x"d1", x"e1", x"c9", x"79", x"0e", x"c1", x"ed", x"79", x"ed", x"41", x"ed", x"59", 
	x"ed", x"51", x"3e", x"00", x"d3", x"c7", x"db", x"c7", x"e6", x"80", x"20", x"fa", x"01", x"c0", x"00", x"ed", 
	x"b2", x"ed", x"b2", x"c9", x"79", x"0e", x"c1", x"ed", x"79", x"ed", x"41", x"ed", x"59", x"ed", x"51", x"3e", 
	x"01", x"d3", x"c7", x"01", x"c0", x"00", x"ed", x"b3", x"ed", x"b3", x"db", x"c7", x"e6", x"80", x"20", x"fa", 
	x"c9", x"dd", x"21", x"f6", x"ff", x"dd", x"39", x"dd", x"71", x"00", x"dd", x"70", x"01", x"e5", x"36", x"06", 
	x"23", x"dd", x"4e", x"00", x"0d", x"0d", x"06", x"00", x"e5", x"d1", x"13", x"36", x"01", x"ed", x"b0", x"36", 
	x"03", x"23", x"e1", x"e5", x"dd", x"5e", x"00", x"16", x"00", x"1d", x"19", x"11", x"20", x"00", x"19", x"dd", 
	x"46", x"01", x"05", x"05", x"36", x"02", x"19", x"10", x"fb", x"e1", x"11", x"20", x"00", x"19", x"dd", x"46", 
	x"01", x"05", x"05", x"36", x"02", x"19", x"10", x"fb", x"36", x"04", x"23", x"dd", x"4e", x"00", x"0d", x"0d", 
	x"06", x"00", x"e5", x"d1", x"13", x"36", x"01", x"ed", x"b0", x"36", x"05", x"23", x"c9", x"21", x"00", x"f0", 
	x"11", x"01", x"f0", x"01", x"ff", x"01", x"36", x"20", x"ed", x"b0", x"c9", x"21", x"00", x"f2", x"11", x"01", 
	x"f2", x"01", x"ff", x"01", x"77", x"ed", x"b0", x"c9", x"7c", x"cd", x"21", x"02", x"7d", x"cd", x"21", x"02", 
	x"c9", x"f5", x"cb", x"3f", x"cb", x"3f", x"cb", x"3f", x"cb", x"3f", x"cd", x"2e", x"02", x"f1", x"e6", x"0f", 
	x"fe", x"0a", x"38", x"05", x"c6", x"37", x"12", x"13", x"c9", x"c6", x"30", x"12", x"13", x"c9", x"2e", x"00", 
	x"55", x"cb", x"24", x"30", x"01", x"6b", x"06", x"07", x"29", x"30", x"01", x"19", x"10", x"fa", x"c9", x"af", 
	x"06", x"10", x"29", x"17", x"b9", x"38", x"02", x"91", x"2c", x"10", x"f7", x"c9", x"c5", x"e5", x"77", x"e5", 
	x"d1", x"13", x"06", x"00", x"0d", x"ed", x"b0", x"e1", x"c1", x"11", x"20", x"00", x"19", x"10", x"ed", x"c9", 
	x"e5", x"c5", x"60", x"59", x"cd", x"3e", x"02", x"29", x"11", x"04", x"00", x"19", x"e5", x"c1", x"cd", x"7e", 
	x"07", x"e5", x"dd", x"e1", x"c1", x"d1", x"dd", x"73", x"00", x"dd", x"72", x"01", x"dd", x"71", x"02", x"dd", 
	x"70", x"03", x"11", x"04", x"00", x"19", x"eb", x"dd", x"4e", x"00", x"dd", x"46", x"01", x"21", x"00", x"f2", 
	x"09", x"cd", x"b5", x"02", x"dd", x"4e", x"00", x"dd", x"46", x"01", x"21", x"00", x"f0", x"09", x"cd", x"b5", 
	x"02", x"dd", x"e5", x"e1", x"c9", x"dd", x"46", x"03", x"c5", x"e5", x"06", x"00", x"dd", x"4e", x"02", x"ed", 
	x"b0", x"e1", x"01", x"20", x"00", x"09", x"c1", x"10", x"ef", x"c9", x"e5", x"dd", x"e1", x"21", x"00", x"f2", 
	x"dd", x"5e", x"00", x"dd", x"56", x"01", x"19", x"eb", x"01", x"04", x"00", x"dd", x"e5", x"e1", x"09", x"cd", 
	x"f9", x"02", x"e5", x"21", x"00", x"f0", x"dd", x"5e", x"00", x"dd", x"56", x"01", x"19", x"eb", x"e1", x"cd", 
	x"f9", x"02", x"dd", x"e5", x"e1", x"cd", x"f1", x"07", x"c9", x"dd", x"46", x"03", x"c5", x"d5", x"06", x"00", 
	x"dd", x"4e", x"02", x"ed", x"b0", x"d1", x"e5", x"21", x"20", x"00", x"19", x"eb", x"e1", x"c1", x"10", x"ec", 
	x"c9", x"7e", x"b7", x"28", x"09", x"12", x"23", x"13", x"0d", x"79", x"b7", x"20", x"f4", x"c9", x"eb", x"78", 
	x"41", x"36", x"20", x"23", x"10", x"fb", x"47", x"c9", x"7e", x"12", x"23", x"13", x"b7", x"20", x"f9", x"c9", 
	x"d5", x"11", x"00", x"00", x"7e", x"b7", x"28", x"09", x"fe", x"2e", x"20", x"02", x"e5", x"d1", x"23", x"18", 
	x"f3", x"eb", x"d1", x"c9", x"c5", x"7e", x"b7", x"28", x"11", x"cd", x"5f", x"03", x"4f", x"1a", x"cd", x"5f", 
	x"03", x"b9", x"20", x"04", x"23", x"13", x"18", x"ed", x"c1", x"c9", x"4f", x"1a", x"b9", x"18", x"f9", x"fe", 
	x"61", x"d8", x"fe", x"7b", x"d0", x"e6", x"5f", x"c9", x"00", x"00", x"19", x"00", x"00", x"00", x"15", x"00", 
	x"13", x"00", x"11", x"00", x"12", x"00", x"1c", x"00", x"00", x"00", x"1a", x"00", x"18", x"00", x"16", x"00", 
	x"14", x"00", x"09", x"00", x"01", x"00", x"00", x"00", x"00", x"00", x"06", x"07", x"02", x"00", x"00", x"00", 
	x"04", x"05", x"51", x"00", x"31", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5a", x"00", x"53", x"00", 
	x"41", x"00", x"57", x"00", x"32", x"00", x"00", x"00", x"00", x"00", x"43", x"00", x"58", x"00", x"44", x"00", 
	x"45", x"00", x"34", x"00", x"33", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"56", x"00", x"46", x"00", 
	x"54", x"00", x"52", x"00", x"35", x"00", x"00", x"00", x"00", x"00", x"4e", x"00", x"42", x"00", x"48", x"00", 
	x"47", x"00", x"59", x"00", x"36", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4d", x"00", x"4a", x"00", 
	x"55", x"00", x"37", x"00", x"38", x"00", x"00", x"00", x"00", x"00", x"0a", x"00", x"4b", x"00", x"49", x"00", 
	x"4f", x"00", x"30", x"00", x"39", x"00", x"00", x"00", x"00", x"00", x"0b", x"00", x"2b", x"5d", x"4c", x"00", 
	x"0e", x"00", x"50", x"00", x"0c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1f", x"00", x"00", x"00", 
	x"1d", x"00", x"0f", x"00", x"00", x"00", x"00", x"00", x"3b", x"00", x"03", x"00", x"0d", x"3c", x"1e", x"00", 
	x"00", x"00", x"3a", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"61", x"26", x"00", x"00", x"64", x"21", 
	x"67", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"29", x"5f", x"2a", x"62", x"24", x"65", x"00", 
	x"66", x"22", x"68", x"23", x"10", x"00", x"00", x"00", x"1b", x"00", x"5e", x"00", x"63", x"27", x"5b", x"00", 
	x"5c", x"00", x"69", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"17", x"00", 
	x"00", x"00", x"60", x"7e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"08", x"08", x"09", x"09", x"2c", x"3c", x"2e", x"3e", x"2d", x"5f", x"0a", x"0a", x"3b", x"3a", x"3d", x"2b", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5b", x"7b", x"5d", x"7d", x"27", x"22", 
	x"20", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"2f", x"3f", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"30", x"29", x"31", x"21", x"32", x"40", x"33", x"23", x"34", x"24", x"35", x"25", x"36", x"5e", x"37", x"26", 
	x"38", x"2a", x"39", x"28", x"5c", x"7c", x"00", x"00", x"0d", x"0d", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"61", x"41", x"62", x"42", x"63", x"43", x"64", x"44", x"65", x"45", x"66", x"46", x"67", x"47", 
	x"68", x"48", x"69", x"49", x"6a", x"4a", x"6b", x"4b", x"6c", x"4c", x"6d", x"4d", x"6e", x"4e", x"6f", x"4f", 
	x"70", x"50", x"71", x"51", x"72", x"52", x"73", x"53", x"74", x"54", x"75", x"55", x"76", x"56", x"77", x"57", 
	x"78", x"58", x"79", x"59", x"7a", x"5a", x"2d", x"2d", x"2a", x"2a", x"2f", x"2f", x"2b", x"2b", x"2e", x"2e", 
	x"30", x"30", x"31", x"31", x"32", x"32", x"33", x"33", x"34", x"34", x"35", x"35", x"36", x"36", x"37", x"37", 
	x"38", x"38", x"39", x"39", x"fd", x"21", x"fc", x"ff", x"fd", x"39", x"fd", x"f9", x"fd", x"6e", x"10", x"fd", 
	x"66", x"11", x"01", x"00", x"00", x"7e", x"b6", x"28", x"05", x"03", x"23", x"23", x"18", x"f7", x"fd", x"71", 
	x"00", x"fd", x"70", x"01", x"af", x"fd", x"77", x"02", x"fd", x"77", x"03", x"fd", x"4e", x"0c", x"fd", x"46", 
	x"0d", x"fd", x"6e", x"0e", x"fd", x"66", x"0f", x"fd", x"7e", x"08", x"11", x"00", x"f2", x"19", x"cd", x"5c", 
	x"02", x"cd", x"80", x"06", x"cd", x"ae", x"06", x"cd", x"e6", x"06", x"cd", x"14", x"07", x"fd", x"7e", x"09", 
	x"cd", x"e7", x"06", x"cd", x"3b", x"01", x"f5", x"fd", x"7e", x"08", x"cd", x"e7", x"06", x"f1", x"fd", x"5e", 
	x"0a", x"fd", x"56", x"0b", x"fe", x"4f", x"20", x"03", x"c3", x"4a", x"06", x"fe", x"23", x"28", x"60", x"fe", 
	x"24", x"28", x"62", x"fe", x"0d", x"20", x"03", x"c3", x"4a", x"06", x"fe", x"10", x"28", x"12", x"fe", x"25", 
	x"28", x"59", x"fe", x"26", x"28", x"5d", x"fe", x"27", x"28", x"65", x"fe", x"28", x"28", x"6d", x"18", x"b1", 
	x"1e", x"ff", x"53", x"c3", x"4a", x"06", x"7a", x"e6", x"80", x"28", x"03", x"11", x"00", x"00", x"fd", x"6e", 
	x"00", x"fd", x"66", x"01", x"b7", x"ed", x"52", x"30", x"07", x"fd", x"5e", x"00", x"fd", x"56", x"01", x"1b", 
	x"fd", x"6e", x"10", x"fd", x"66", x"11", x"19", x"19", x"d5", x"5e", x"23", x"56", x"eb", x"d1", x"7e", x"fe", 
	x"2d", x"20", x"03", x"eb", x"09", x"eb", x"fd", x"73", x"0a", x"fd", x"72", x"0b", x"c3", x"81", x"05", x"1b", 
	x"01", x"ff", x"ff", x"18", x"c1", x"13", x"01", x"01", x"00", x"18", x"bb", x"11", x"00", x"00", x"01", x"01", 
	x"00", x"18", x"b3", x"fd", x"5e", x"00", x"fd", x"56", x"01", x"1b", x"01", x"ff", x"ff", x"18", x"a7", x"fd", 
	x"6e", x"0d", x"26", x"00", x"19", x"eb", x"01", x"01", x"00", x"18", x"9b", x"fd", x"6e", x"0d", x"26", x"00", 
	x"eb", x"b7", x"ed", x"52", x"eb", x"01", x"ff", x"ff", x"18", x"8c", x"fd", x"6e", x"06", x"fd", x"66", x"07", 
	x"7d", x"b4", x"28", x"21", x"e5", x"dd", x"e1", x"7a", x"e6", x"80", x"28", x"05", x"21", x"00", x"00", x"18", 
	x"08", x"fd", x"6e", x"10", x"fd", x"66", x"11", x"19", x"19", x"fd", x"e5", x"cd", x"7e", x"06", x"fd", x"e1", 
	x"28", x"03", x"c3", x"81", x"05", x"fd", x"21", x"04", x"00", x"fd", x"39", x"fd", x"f9", x"c9", x"dd", x"e9", 
	x"fd", x"6e", x"0a", x"fd", x"66", x"0b", x"7c", x"e6", x"80", x"28", x"09", x"fd", x"36", x"0a", x"00", x"fd", 
	x"36", x"0b", x"00", x"c9", x"eb", x"fd", x"6e", x"00", x"fd", x"66", x"01", x"2b", x"b7", x"ed", x"52", x"d0", 
	x"fd", x"6e", x"00", x"fd", x"66", x"01", x"2b", x"fd", x"75", x"0a", x"fd", x"74", x"0b", x"c9", x"fd", x"6e", 
	x"0a", x"fd", x"66", x"0b", x"fd", x"5e", x"02", x"fd", x"56", x"03", x"e5", x"d5", x"b7", x"ed", x"52", x"d1", 
	x"e1", x"30", x"07", x"fd", x"75", x"02", x"fd", x"74", x"03", x"c9", x"fd", x"4e", x"0d", x"06", x"00", x"0d", 
	x"eb", x"09", x"eb", x"b7", x"ed", x"52", x"d8", x"c8", x"fd", x"5e", x"02", x"fd", x"56", x"03", x"19", x"fd", 
	x"75", x"02", x"fd", x"74", x"03", x"c9", x"c9", x"fd", x"6e", x"0a", x"fd", x"66", x"0b", x"fd", x"5e", x"02", 
	x"fd", x"56", x"03", x"b7", x"ed", x"52", x"5d", x"26", x"20", x"cd", x"3e", x"02", x"11", x"00", x"f2", x"19", 
	x"fd", x"5e", x"0e", x"fd", x"56", x"0f", x"19", x"e5", x"d1", x"13", x"06", x"00", x"fd", x"4e", x"0c", x"0d", 
	x"77", x"ed", x"b0", x"c9", x"21", x"00", x"f0", x"fd", x"5e", x"0e", x"fd", x"56", x"0f", x"19", x"eb", x"fd", 
	x"6e", x"10", x"fd", x"66", x"11", x"fd", x"4e", x"02", x"fd", x"46", x"03", x"09", x"09", x"e5", x"dd", x"e1", 
	x"fd", x"46", x"0d", x"dd", x"6e", x"00", x"dd", x"66", x"01", x"7d", x"b4", x"28", x"18", x"7e", x"fe", x"2d", 
	x"20", x"1a", x"d5", x"d5", x"e1", x"13", x"c5", x"fd", x"4e", x"0c", x"0d", x"06", x"00", x"36", x"01", x"ed", 
	x"b0", x"c1", x"d1", x"18", x"0f", x"21", x"70", x"07", x"dd", x"2b", x"dd", x"2b", x"d5", x"fd", x"4e", x"0c", 
	x"cd", x"11", x"03", x"d1", x"21", x"20", x"00", x"19", x"eb", x"dd", x"23", x"dd", x"23", x"10", x"c4", x"c9", 
	x"00", x"21", x"00", x"00", x"22", x"00", x"42", x"21", x"e2", x"42", x"22", x"02", x"42", x"c9", x"dd", x"21", 
	x"00", x"00", x"dd", x"39", x"3e", x"00", x"b0", x"20", x"07", x"79", x"fe", x"02", x"30", x"02", x"0e", x"02", 
	x"dd", x"36", x"f6", x"00", x"dd", x"36", x"f7", x"00", x"2a", x"00", x"42", x"7c", x"b5", x"28", x"31", x"5e", 
	x"23", x"56", x"23", x"7b", x"91", x"7a", x"98", x"30", x"0d", x"dd", x"75", x"f6", x"dd", x"74", x"f7", x"5e", 
	x"23", x"56", x"23", x"eb", x"18", x"e5", x"e5", x"5e", x"23", x"56", x"23", x"dd", x"6e", x"f6", x"dd", x"66", 
	x"f7", x"7d", x"b4", x"28", x"05", x"73", x"23", x"72", x"18", x"04", x"eb", x"22", x"00", x"42", x"e1", x"c9", 
	x"2a", x"02", x"42", x"09", x"23", x"23", x"11", x"e2", x"7a", x"7b", x"95", x"7a", x"9c", x"38", x"0e", x"2a", 
	x"02", x"42", x"71", x"23", x"70", x"23", x"e5", x"09", x"22", x"02", x"42", x"e1", x"c9", x"21", x"00", x"00", 
	x"c9", x"2b", x"46", x"2b", x"4e", x"e5", x"09", x"23", x"23", x"eb", x"2a", x"02", x"42", x"7a", x"bc", x"20", 
	x"09", x"7b", x"bd", x"20", x"05", x"e1", x"22", x"02", x"42", x"c9", x"e1", x"ed", x"5b", x"00", x"42", x"22", 
	x"00", x"42", x"23", x"23", x"73", x"23", x"72", x"c9", x"3c", x"65", x"6a", x"65", x"63", x"74", x"3e", x"00", 
	x"fd", x"21", x"f4", x"ff", x"fd", x"39", x"fd", x"f9", x"fd", x"77", x"00", x"fd", x"73", x"06", x"fd", x"72", 
	x"07", x"3e", x"ff", x"fd", x"77", x"02", x"fd", x"77", x"03", x"7c", x"e6", x"80", x"20", x"0e", x"29", x"29", 
	x"29", x"29", x"29", x"eb", x"2a", x"26", x"42", x"19", x"11", x"0a", x"00", x"19", x"fd", x"75", x"04", x"fd", 
	x"74", x"05", x"21", x"42", x"00", x"01", x"1c", x"0c", x"cd", x"70", x"02", x"fd", x"75", x"08", x"fd", x"74", 
	x"09", x"21", x"42", x"f2", x"01", x"1c", x"0c", x"3e", x"cf", x"cd", x"5c", x"02", x"21", x"42", x"f0", x"01", 
	x"1c", x"0c", x"cd", x"a1", x"01", x"2a", x"28", x"42", x"29", x"23", x"23", x"23", x"23", x"e5", x"c1", x"cd", 
	x"7e", x"07", x"fd", x"75", x"0a", x"fd", x"74", x"0b", x"e5", x"dd", x"e1", x"fd", x"7e", x"00", x"b7", x"28", 
	x"0d", x"21", x"18", x"08", x"dd", x"75", x"00", x"dd", x"74", x"01", x"dd", x"23", x"dd", x"23", x"2a", x"26", 
	x"42", x"11", x"0a", x"00", x"19", x"ed", x"4b", x"28", x"42", x"7e", x"b7", x"28", x"3b", x"fd", x"5e", x"06", 
	x"fd", x"56", x"07", x"e5", x"cd", x"84", x"09", x"e1", x"20", x"2e", x"fd", x"7e", x"04", x"bd", x"20", x"1e", 
	x"fd", x"7e", x"05", x"bc", x"20", x"18", x"e5", x"dd", x"e5", x"e1", x"fd", x"5e", x"0a", x"fd", x"56", x"0b", 
	x"b7", x"ed", x"52", x"cb", x"3c", x"cb", x"1d", x"fd", x"75", x"02", x"fd", x"74", x"03", x"e1", x"dd", x"75", 
	x"00", x"dd", x"74", x"01", x"dd", x"23", x"dd", x"23", x"11", x"20", x"00", x"19", x"0b", x"78", x"b1", x"20", 
	x"b8", x"af", x"dd", x"77", x"00", x"dd", x"77", x"01", x"fd", x"e5", x"fd", x"6e", x"0a", x"fd", x"66", x"0b", 
	x"e5", x"21", x"63", x"00", x"e5", x"21", x"1a", x"0a", x"e5", x"fd", x"6e", x"02", x"fd", x"66", x"03", x"e5", 
	x"21", x"cf", x"b0", x"e5", x"21", x"00", x"00", x"e5", x"cd", x"44", x"05", x"fd", x"21", x"0c", x"00", x"fd", 
	x"39", x"fd", x"f9", x"fd", x"e1", x"7a", x"e6", x"80", x"20", x"3d", x"fd", x"7e", x"00", x"b7", x"28", x"04", 
	x"7a", x"b3", x"28", x"30", x"fd", x"6e", x"0a", x"fd", x"66", x"0b", x"19", x"19", x"5e", x"23", x"56", x"eb", 
	x"11", x"0a", x"00", x"b7", x"ed", x"52", x"ed", x"5b", x"26", x"42", x"b7", x"ed", x"52", x"cb", x"3c", x"cb", 
	x"1d", x"cb", x"3c", x"cb", x"1d", x"cb", x"3c", x"cb", x"1d", x"cb", x"3c", x"cb", x"1d", x"cb", x"3c", x"cb", 
	x"1d", x"eb", x"18", x"03", x"11", x"fe", x"ff", x"d5", x"fd", x"6e", x"0a", x"fd", x"66", x"0b", x"cd", x"f1", 
	x"07", x"fd", x"6e", x"08", x"fd", x"66", x"09", x"cd", x"ca", x"02", x"d1", x"fd", x"21", x"0c", x"00", x"fd", 
	x"39", x"fd", x"f9", x"c9", x"7a", x"b3", x"c8", x"cd", x"30", x"03", x"7c", x"b5", x"20", x"03", x"f6", x"01", 
	x"c9", x"23", x"e5", x"cd", x"44", x"03", x"e1", x"c8", x"1a", x"b7", x"13", x"20", x"fb", x"1a", x"b7", x"20", 
	x"f1", x"f6", x"01", x"c9", x"46", x"50", x"47", x"41", x"42", x"65", x"65", x"20", x"76", x"32", x"2e", x"30", 
	x"2e", x"31", x"2a", x"42", x"4a", x"42", x"6a", x"42", x"fa", x"09", x"fc", x"09", x"00", x"00", x"64", x"73", 
	x"34", x"30", x"00", x"73", x"73", x"38", x"30", x"00", x"64", x"73", x"38", x"30", x"00", x"64", x"73", x"38", 
	x"32", x"00", x"64", x"73", x"38", x"34", x"00", x"64", x"73", x"38", x"42", x"00", x"68", x"64", x"30", x"00", 
	x"00", x"68", x"64", x"31", x"00", x"00", x"48", x"44", x"31", x"3a", x"00", x"46", x"44", x"30", x"3a", x"00", 
	x"46", x"44", x"31", x"3a", x"00", x"46", x"44", x"32", x"3a", x"00", x"2d", x"00", x"52", x"65", x"73", x"65", 
	x"74", x"00", x"31", x"00", x"80", x"cd", x"71", x"07", x"3e", x"00", x"cd", x"0b", x"02", x"cd", x"fd", x"01", 
	x"db", x"c7", x"e6", x"40", x"20", x"fa", x"cd", x"58", x"0b", x"cd", x"88", x"0b", x"cd", x"4a", x"0c", x"cd", 
	x"ba", x"0c", x"21", x"e6", x"09", x"11", x"2a", x"42", x"ed", x"4b", x"1a", x"42", x"cd", x"de", x"0b", x"21", 
	x"eb", x"09", x"11", x"4a", x"42", x"ed", x"4b", x"1e", x"42", x"cd", x"de", x"0b", x"21", x"f0", x"09", x"11", 
	x"6a", x"42", x"ed", x"4b", x"20", x"42", x"cd", x"de", x"0b", x"21", x"00", x"f2", x"01", x"20", x"07", x"3e", 
	x"cf", x"cd", x"5c", x"02", x"21", x"00", x"f0", x"01", x"20", x"07", x"cd", x"a1", x"01", x"21", x"a4", x"09", 
	x"11", x"09", x"f0", x"01", x"0e", x"00", x"ed", x"b0", x"21", x"b2", x"09", x"e5", x"21", x"21", x"00", x"e5", 
	x"21", x"1e", x"05", x"e5", x"21", x"00", x"00", x"e5", x"21", x"cf", x"b0", x"e5", x"21", x"8e", x"0a", x"e5", 
	x"cd", x"44", x"05", x"18", x"fe", x"7e", x"cd", x"21", x"02", x"23", x"13", x"10", x"f8", x"c9", x"7a", x"e6", 
	x"80", x"20", x"1d", x"7b", x"fe", x"00", x"28", x"1f", x"fe", x"01", x"28", x"2d", x"fe", x"02", x"28", x"3b", 
	x"fe", x"04", x"28", x"03", x"f6", x"01", x"c9", x"3e", x"00", x"d3", x"81", x"d3", x"ff", x"f6", x"01", x"c9", 
	x"3e", x"00", x"d3", x"81", x"f6", x"01", x"c9", x"2a", x"1a", x"42", x"11", x"30", x"0b", x"3e", x"01", x"cd", 
	x"20", x"08", x"21", x"2f", x"42", x"0e", x"01", x"18", x"24", x"2a", x"1e", x"42", x"11", x"39", x"0b", x"3e", 
	x"01", x"cd", x"20", x"08", x"21", x"4f", x"42", x"0e", x"03", x"18", x"12", x"2a", x"20", x"42", x"11", x"39", 
	x"0b", x"3e", x"01", x"cd", x"20", x"08", x"21", x"6f", x"42", x"0e", x"04", x"18", x"00", x"7a", x"e6", x"80", 
	x"28", x"12", x"7b", x"fe", x"fe", x"28", x"03", x"f6", x"01", x"c9", x"36", x"2d", x"23", x"36", x"00", x"11", 
	x"ff", x"ff", x"18", x"16", x"d5", x"e5", x"eb", x"29", x"29", x"29", x"29", x"29", x"ed", x"5b", x"26", x"42", 
	x"19", x"11", x"0a", x"00", x"19", x"d1", x"cd", x"28", x"03", x"d1", x"c5", x"21", x"18", x"42", x"06", x"00", 
	x"09", x"09", x"73", x"23", x"72", x"c1", x"79", x"cd", x"06", x"0c", x"cd", x"70", x"0b", x"f6", x"01", x"c9", 
	x"68", x"64", x"30", x"00", x"68", x"64", x"31", x"00", x"00", x"64", x"73", x"34", x"30", x"00", x"73", x"73", 
	x"38", x"30", x"00", x"64", x"73", x"38", x"30", x"00", x"64", x"73", x"38", x"32", x"00", x"64", x"73", x"38", 
	x"34", x"00", x"64", x"73", x"38", x"62", x"00", x"00", x"11", x"00", x"00", x"01", x"00", x"00", x"21", x"00", 
	x"40", x"cd", x"67", x"01", x"21", x"00", x"40", x"11", x"04", x"42", x"01", x"22", x"00", x"ed", x"b0", x"c9", 
	x"21", x"04", x"42", x"11", x"00", x"40", x"01", x"22", x"00", x"ed", x"b0", x"11", x"00", x"00", x"01", x"00", 
	x"00", x"21", x"00", x"40", x"cd", x"84", x"01", x"c9", x"3a", x"0e", x"42", x"cb", x"27", x"47", x"0e", x"00", 
	x"cd", x"7e", x"07", x"22", x"26", x"42", x"ed", x"4b", x"0a", x"42", x"ed", x"5b", x"0c", x"42", x"3a", x"0e", 
	x"42", x"f5", x"c5", x"d5", x"cd", x"67", x"01", x"d1", x"c1", x"e5", x"21", x"01", x"00", x"09", x"e5", x"c1", 
	x"21", x"00", x"00", x"ed", x"5a", x"eb", x"e1", x"f1", x"d6", x"01", x"20", x"e5", x"dd", x"2a", x"26", x"42", 
	x"01", x"00", x"00", x"11", x"20", x"00", x"dd", x"7e", x"00", x"dd", x"b6", x"01", x"dd", x"b6", x"02", x"dd", 
	x"b6", x"03", x"28", x"05", x"dd", x"19", x"03", x"18", x"ed", x"ed", x"43", x"28", x"42", x"c9", x"cd", x"28", 
	x"03", x"eb", x"2b", x"36", x"20", x"23", x"78", x"e6", x"80", x"28", x"06", x"36", x"2d", x"23", x"36", x"00", 
	x"c9", x"eb", x"c5", x"e1", x"29", x"29", x"29", x"29", x"29", x"01", x"0a", x"00", x"09", x"ed", x"4b", x"26", 
	x"42", x"09", x"cd", x"28", x"03", x"c9", x"e5", x"c5", x"f5", x"7a", x"e6", x"80", x"28", x"0e", x"3e", x"00", 
	x"d3", x"c1", x"d3", x"c1", x"d3", x"c1", x"d3", x"c1", x"3e", x"08", x"18", x"19", x"eb", x"29", x"29", x"29", 
	x"29", x"29", x"ed", x"5b", x"26", x"42", x"19", x"e5", x"01", x"c1", x"04", x"ed", x"b3", x"e1", x"11", x"0a", 
	x"00", x"19", x"cd", x"d0", x"0c", x"cb", x"27", x"cb", x"27", x"cb", x"27", x"47", x"f1", x"fe", x"03", x"38", 
	x"01", x"3c", x"f6", x"80", x"b0", x"d3", x"c7", x"c1", x"e1", x"c9", x"21", x"18", x"42", x"06", x"07", x"5e", 
	x"23", x"56", x"23", x"3e", x"07", x"90", x"cd", x"06", x"0c", x"10", x"f4", x"c9", x"f6", x"80", x"d3", x"d0", 
	x"d5", x"21", x"00", x"80", x"11", x"01", x"80", x"01", x"ff", x"3f", x"36", x"00", x"ed", x"b0", x"d1", x"7a", 
	x"e6", x"80", x"20", x"42", x"eb", x"29", x"29", x"29", x"29", x"29", x"ed", x"5b", x"26", x"42", x"19", x"11", 
	x"aa", x"42", x"01", x"04", x"00", x"ed", x"b0", x"7e", x"3d", x"e6", x"1f", x"3c", x"47", x"21", x"00", x"80", 
	x"c5", x"ed", x"4b", x"aa", x"42", x"ed", x"5b", x"ac", x"42", x"cd", x"67", x"01", x"eb", x"2a", x"aa", x"42", 
	x"01", x"01", x"00", x"09", x"22", x"aa", x"42", x"2a", x"ac", x"42", x"01", x"00", x"00", x"ed", x"4a", x"22", 
	x"ac", x"42", x"eb", x"c1", x"10", x"da", x"af", x"d3", x"d0", x"c9", x"21", x"12", x"42", x"06", x"03", x"5e", 
	x"23", x"56", x"23", x"3e", x"03", x"90", x"c5", x"e5", x"cd", x"5c", x"0c", x"e1", x"c1", x"10", x"f0", x"c9", 
	x"cd", x"30", x"03", x"7c", x"b5", x"20", x"03", x"3e", x"08", x"c9", x"23", x"06", x"08", x"11", x"be", x"09", 
	x"eb", x"e5", x"d5", x"cd", x"44", x"03", x"d1", x"e1", x"28", x"08", x"c5", x"01", x"05", x"00", x"09", x"c1", 
	x"10", x"ef", x"3e", x"08", x"90", x"c9", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"
	
	);
begin

	process (clock)
	begin
		if rising_edge(clock) then
			if clken='1' then
				dout <= rom(to_integer(unsigned(addr)));
			end if;
		end if;
	end process;
end;

